library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

-- clock division factor: 125
-- signal frequency division factor: 250
-- depth: 6 periods
entity lpf_rom_125_250 is
	port(addr1,addr2: in unsigned(6 downto 0);
			clk: in std_logic;
			--output consists of 12 8-bit signed 2's complement
			--fractions (all bits fractional);
			--data[0] is sinc(0)&sinc(1)&sinc(2)...
			--data[1] is sinc(0+1/125)&sinc(1+1/125)&...
			q1,q2: out signed(95 downto 0));
end entity;
architecture a of lpf_rom_125_250 is
	type rom1t is array(0 to 124) of signed(95 downto 0);
	signal rom1: rom1t := (
X"f9000900f4001000e500517f",
X"f9000900f4001000e5ff507f",
X"f9000900f4001001e5ff507f",
X"f9000900f4ff1001e5fe4f7f",
X"f9000901f5ff1001e5fe4e7f",
X"f9ff0901f5ff1001e5fe4e7f",
X"f9ff0901f5ff1002e6fd4d7f",
X"f9ff0901f5ff1002e6fd4c7f",
X"f9ff0901f5ff1002e6fc4c7f",
X"f9ff0901f5fe1002e6fc4b7f",
X"f9ff0901f5fe1002e6fb4a7f",
X"f9ff0901f5fe1003e6fb4a7f",
X"f9ff0902f5fe1003e6fa497f",
X"f9ff0902f5fe1003e6fa487e",
X"f9ff0902f5fe1003e6f9487e",
X"f9ff0902f5fe1004e7f9477e",
X"f9fe0902f5fd0f04e7f8467e",
X"f9fe0902f5fd0f04e7f8467e",
X"f9fe0902f5fd0f04e7f8457e",
X"f9fe0902f5fd0f05e7f7447e",
X"f9fe0902f5fd0f05e7f7447e",
X"f9fe0903f5fd0f05e7f6437e",
X"f9fe0803f5fc0f05e8f6427d",
X"f9fe0803f5fc0f06e8f5417d",
X"f9fe0803f5fc0f06e8f5417d",
X"f9fe0803f5fc0f06e8f5407d",
X"f9fd0803f5fc0f06e8f43f7d",
X"f9fd0803f5fc0f06e8f43f7d",
X"f9fd0803f5fc0f07e8f33e7c",
X"f9fd0804f6fb0e07e9f33d7c",
X"f9fd0804f6fb0e07e9f33d7c",
X"f9fd0804f6fb0e07e9f23c7c",
X"f9fd0804f6fb0e07e9f23b7c",
X"f9fd0804f6fb0e08e9f23b7b",
X"f9fd0804f6fb0e08eaf13a7b",
X"fafd0804f6fb0e08eaf1397b",
X"fafd0804f6fa0e08eaf1387b",
X"fafc0804f6fa0e08eaf0387a",
X"fafc0804f6fa0e09eaf0377a",
X"fafc0805f6fa0d09eaf0367a",
X"fafc0805f6fa0d09ebef367a",
X"fafc0805f6fa0d09ebef3579",
X"fafc0705f6fa0d09ebef3479",
X"fafc0705f7f90d0aebee3479",
X"fafc0705f7f90d0aebee3379",
X"fafc0705f7f90d0aecee3278",
X"fafc0705f7f90d0aeced3178",
X"fafc0705f7f90c0aeced3178",
X"fafc0705f7f90c0aeced3077",
X"fafc0706f7f90c0bedec2f77",
X"fafb0706f7f90c0bedec2f77",
X"fafb0706f7f80c0bedec2e76",
X"fafb0706f7f80c0bedec2d76",
X"fafb0706f7f80c0bedeb2d76",
X"fafb0706f8f80c0beeeb2c75",
X"fbfb0706f8f80b0ceeeb2b75",
X"fbfb0706f8f80b0ceeeb2b75",
X"fbfb0606f8f80b0ceeea2a74",
X"fbfb0606f8f80b0cefea2974",
X"fbfb0606f8f80b0cefea2974",
X"fbfb0607f8f70b0cefea2873",
X"fbfb0607f8f70b0cefe92773",
X"fbfb0607f8f70a0df0e92673",
X"fbfb0607f8f70a0df0e92672",
X"fbfa0607f9f70a0df0e92572",
X"fbfa0607f9f70a0df0e92471",
X"fbfa0607f9f70a0df1e82471",
X"fbfa0607f9f70a0df1e82371",
X"fbfa0607f9f70a0df1e82270",
X"fbfa0507f9f7090ef1e82270",
X"fcfa0507f9f7090ef2e8216f",
X"fcfa0507f9f6090ef2e7206f",
X"fcfa0507f9f6090ef2e7206e",
X"fcfa0507faf6090ef2e71f6e",
X"fcfa0508faf6090ef3e71e6d",
X"fcfa0508faf6080ef3e71e6d",
X"fcfa0508faf6080ef3e71d6d",
X"fcfa0508faf6080ef3e71c6c",
X"fcfa0508faf6080ff4e61c6c",
X"fcfa0508faf6080ff4e61b6b",
X"fcfa0408faf6080ff4e61a6b",
X"fcfa0408faf6080ff4e61a6a",
X"fcf90408fbf6070ff5e6196a",
X"fdf90408fbf6070ff5e61869",
X"fdf90408fbf5070ff5e61869",
X"fdf90408fbf5070ff5e61768",
X"fdf90408fbf5070ff6e51768",
X"fdf90408fbf5070ff6e51667",
X"fdf90408fbf5060ff6e51567",
X"fdf90408fbf5060ff6e51566",
X"fdf90408fcf5060ff7e51466",
X"fdf90308fcf50610f7e51365",
X"fdf90308fcf50610f7e51365",
X"fdf90309fcf50610f8e51264",
X"fdf90309fcf50510f8e51263",
X"fdf90309fcf50510f8e51163",
X"fef90309fcf50510f8e51062",
X"fef90309fcf50510f9e51062",
X"fef90309fdf50510f9e50f61",
X"fef90309fdf50410f9e50e61",
X"fef90309fdf50410f9e50e60",
X"fef90209fdf50410fae50d60",
X"fef90209fdf50410fae40d5f",
X"fef90209fdf50410fae40c5e",
X"fef90209fdf50410fae40c5e",
X"fef90209fdf50310fbe40b5d",
X"fef90209fef50310fbe40a5d",
X"fef90209fef50310fbe40a5c",
X"fff90209fef40310fce4095b",
X"fff90209fef40310fce4095b",
X"fff90209fef40310fce4085a",
X"fff90109fef40210fce4075a",
X"fff90109fef40210fde40759",
X"fff90109fef40210fde40658",
X"fff90109fff40210fde50658",
X"fff90109fff40210fde50557",
X"fff90109fff40210fee50557",
X"fff90109fff40110fee50456",
X"fff90109fff40110fee50455",
X"fff90109fff40110fee50355",
X"00f90109fff40110ffe50354",
X"00f90009fff40110ffe50253",
X"00f9000900f40110ffe50253",
X"00f9000900f40010ffe50152",
X"00f9000900f4001000e50151"
);
	signal addr11,addr21: unsigned(6 downto 0);
begin
	addr11 <= addr1 when rising_edge(clk);
	addr21 <= addr2 when rising_edge(clk);
	q1 <= rom1(to_integer(addr11)) when rising_edge(clk);
	q2 <= rom1(to_integer(addr21)) when rising_edge(clk);
end architecture;
