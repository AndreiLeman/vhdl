altlvds_tx1_inst : altlvds_tx1 PORT MAP (
		tx_in	 => tx_in_sig,
		tx_inclock	 => tx_inclock_sig,
		tx_out	 => tx_out_sig
	);
