library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
entity sinc_rom is
	port(addr1,addr2: in unsigned(7 downto 0);
			clk1,clk2: in std_logic;
			--output consists of 6 24-bit signed 2's complement
			--fractions (all bits fractional);
			--data[0] is sinc(0)&sinc(1)&sinc(2)...
			--data[1] is sinc(0+1/192)&sinc(1+1/192)&...
			q1,q2: out signed(143 downto 0));
end entity;
architecture a of sinc_rom is
	type rom1t is array(0 to 255) of signed(143 downto 0);
	signal rom1: rom1t := (
X"7fffcbffc020001ff8ffeaae000ffefff335",
X"7ffe26ff4121005fb7ffc021002fedffd9a6",
X"7ffadcfec325009f33ff95b2004fcbffc023",
X"7ff5edfe462e00de69ff6b64006f96ffa6ac",
X"7fef59fdca3d011d59ff4137008f4cff8d43",
X"7fe720fd4f54015bffff172e00aeedff73e9",
X"7fdd43fcd576019a59feed4900ce78ff5a9e",
X"7fd1c1fc5ca401d867fec38b00edebff4163",
X"7fc49cfbe4df021625fe99f4010d46ff283a",
X"7fb5d3fb6e2a025393fe7087012c86ff0f23",
X"7fa566faf8860290adfe4744014bacfef620",
X"7f9356fa83f402cd72fe1e2d016ab5fedd30",
X"7f7fa4fa10770309e0fdf5440189a1fec456",
X"7f6a50f99e0f0345f5fdcc8901a86efeab92",
X"7f535af92cbf0381b0fda3ff01c71cfe92e4",
X"7f3ac2f8bc8703bd0efd7ba701e5aafe7a4f",
X"7f208bf84d6a03f80efd5382020415fe61d2",
X"7f04b3f7df680432aefd2b9102225efe496f",
X"7ee73cf77284046cebfd03d6024083fe3126",
X"7ec827f706be04a6c5fcdc53025e83fe18f8",
X"7ea773f69c1704e03afcb508027c5dfe00e7",
X"7e8523f63292051947fc8df7029a10fde8f3",
X"7e6136f5ca300551ecfc672102b79afdd11e",
X"7e3badf562f0058a26fc408802d4fbfdb967",
X"7e148af4fcd605c1f4fc1a2d02f232fda1cf",
X"7debcef497e205f954fbf411030f3efd8a59",
X"7dc178f43415063044fbce36032c1dfd7303",
X"7d958bf3d1700666c3fba89c0348d0fd5bd1",
X"7d6806f36ff5069cd0fb8345036553fd44c1",
X"7d38ecf30fa306d268fb5e320381a8fd2dd5",
X"7d083ef2b07e07078bfb3965039dccfd170e",
X"7cd5fcf25284073c36fb14de03b9befd006c",
X"7ca227f1f5b8077068faf09f03d57ffce9f1",
X"7c6cc1f19a1a07a421faccaa03f10cfcd39e",
X"7c35ccf13fab07d75dfaa8fe040c65fcbd72",
X"7bfd47f0e66d080a1cfa859e042789fca76f",
X"7bc335f08e5e083c5dfa628a044277fc9195",
X"7b8797f03782086e1efa3fc4045d2efc7be6",
X"7b4a6fefe1d7089f5dfa1d4d0477adfc6662",
X"7b0bbdef8d6008d01af9fb250491f3fc5109",
X"7acb83ef3a1c090053f9d94f04abfffc3bde",
X"7a89c3eee80d093006f9b7cb04c5d1fc26e0",
X"7a467eee9732095f33f9969904df67fc120f",
X"7a01b6ee478d098dd8f975bc04f8c1fbfd6e",
X"79bb6cedf91e09bbf4f955340511defbe8fc",
X"7973a2edabe509e986f93502052abdfbd4ba",
X"792a5aed5fe40a168cf9152805435dfbc0aa",
X"78df95ed151a0a4306f8f5a5055bbefbacca",
X"789355eccb870a6ef2f8d67c0573defb991e",
X"78459bec832d0a9a50f8b7ad058bbcfb85a4",
X"77f66aec3c0c0ac51df8993905a359fb725e",
X"77a5c4ebf6230aef59f87b2105bab2fb5f4c",
X"7753a9ebb1740b1904f85d6505d1c9fb4c6f",
X"77001deb6dfd0b421bf8400805e89afb39c8",
X"76ab20eb2bc10b6a9ef8230905ff27fb2757",
X"7654b6eaeabe0b928cf8066a06156efb151d",
X"75fcdfeaaaf60bb9e4f7ea2b062b6efb031a",
X"75a39fea6c670be0a5f7ce4e064127faf14f",
X"7548f6ea2f120c06cff7b2d2065699fadfbd",
X"74ece7e9f2f80c2c60f797ba066bc1face65",
X"748f75e9b8170c5157f77d040680a0fabd46",
X"7430a0e97e710c75b4f762b4069536faac62",
X"73d06de946050c9976f748c806a980fa9bb8",
X"736edce90ed30cbc9bf72f4306bd80fa8b4a",
X"730befe8d8db0cdf25f7162306d133fa7b19",
X"72a7aae8a41d0d0110f6fd6c06e49afa6b23",
X"72420ee870980d225ef6e51c06f7b4fa5b6b",
X"71db1fe83e4c0d430cf6cd35070a80fa4bf1",
X"7172dde80d3a0d631cf6b5b7071cfefa3cb4",
X"71094be7dd600d828bf69ea3072f2efa2db7",
X"709e6de7aebf0da159f687fa07410efa1ef8",
X"703244e781560dbf86f671bb07529efa1079",
X"6fc4d2e755250ddd11f65be90763ddfa023a",
X"6f561be72a2c0df9faf646830774ccf9f43b",
X"6ee621e700690e1640f6318a078569f9e67e",
X"6e74e6e6d7dd0e31e2f61cfe0795b5f9d901",
X"6e026de6b0860e4ce0f608e007a5aef9cbc7",
X"6d8eb9e68a650e673af5f53007b554f9bece",
X"6d19cce665790e80f0f5e1f007c4a7f9b219",
X"6ca3a8e641c20e9a00f5cf1e07d3a6f9a5a6",
X"6c2c51e61f3e0eb26bf5bcbd07e251f99976",
X"6bb3c9e5fded0eca2ff5aacc07f0a8f98d8a",
X"6b3a14e5ddce0ee14ef5994b07fea9f981e3",
X"6abf32e5bee10ef7c6f5883c080c56f9767f",
X"6a4329e5a1240f0d97f5779e0819acf96b61",
X"69c5f9e584980f22c2f567720826adf96087",
X"6947a7e5693b0f3745f557b7083357f955f3",
X"68c835e54f0d0f4b20f54870083fabf94ba5",
X"6847a6e5360c0f5e54f5399b084ba7f9419c",
X"67c5fce51e380f70e1f52b3908574df937da",
X"67433be5078f0f82c5f51d4b08629af92e5e",
X"66bf66e4f2120f9401f50fd0086d90f92529",
X"663a7fe4ddbe0fa495f502c908782ef91c3c",
X"65b48ae4ca930fb482f4f636088273f91395",
X"652d89e4b8900fc3c5f4ea18088c5ff90b36",
X"64a581e4a7b30fd261f4de6e0895f3f9031f",
X"641c72e497fc0fe055f4d338089f2ef8fb4f",
X"639262e4896a0feda0f4c87708a810f8f3c8",
X"630753e47bfb0ffa43f4be2c08b098f8ec89",
X"627b47e46fae10063ef4b45508b8c6f8e592",
X"61ee43e46482101192f4aaf308c09bf8dee4",
X"616049e45a75101c3df4a20708c816f8d87f",
X"60d15de45187102641f4999008cf37f8d263",
X"604181e449b7102f9ef4918e08d5fef8cc90",
X"5fb0bae44302103853f48a0208dc6bf8c706",
X"5f1f09e43d68104061f482eb08e27df8c1c5",
X"5e8c73e438e61047c8f47c4a08e835f8bcce",
X"5df8fbe4357d104e89f4761e08ed93f8b820",
X"5d64a3e4332a1054a4f4706708f296f8b3bc",
X"5ccf70e431eb105a18f46b2608f73ef8afa1",
X"5c3965e431c0105ee8f4665908fb8cf8abd0",
X"5ba284e432a8106311f4620208ff80f8a849",
X"5b0ad2e4349f106696f45e21090319f8a50b",
X"5a7251e437a5106976f45ab3090658f8a217",
X"59d906e43bb9106bb3f457bb09093cf89f6d",
X"593ef3e440d8106d4bf45538090bc6f89d0c",
X"58a41ce44701106e41f45329090df5f89af6",
X"580884e44e33106e94f4518e090fcaf89929",
X"576c2fe4566c106e44f45067091145f897a5",
X"56cf20e45fa9106d53f44fb4091266f8966c",
X"56315be469ea106bc1f44f7509132df8957b",
X"5592e2e4752d10698ff44fa909139af894d5",
X"54f3bbe4816f1066bcf450500913aef89477",
X"5453e8e48eb010634af4516a091367f89463",
X"53b36ce49ced105f39f452f70912c8f89498",
X"53124ce4ac24105a8bf454f60911cff89517",
X"52708be4bc5410553ff4576609107ef895de",
X"51ce2be4cd7b104f56f45a49090ed3f896ee",
X"512b32e4df961048d1f45d9c090cd0f89847",
X"5087a2e4f2a51041b1f46160090a75f899e8",
X"4fe37fe506a51039f6f465950907c1f89bd2",
X"4f3ecde51b941031a2f46a3a0904b6f89e04",
X"4e998fe5316f1028b4f46f4e090153f8a07e",
X"4df3c8e54837101f2ff474d108fd99f8a33f",
X"4d4d7ee55fe7101512f47ac308f987f8a649",
X"4ca6b2e5787e100a5ff4812408f51ff8a99a",
X"4bff69e591fb0fff16f487f108f061f8ad32",
X"4b57a6e5ac5a0ff338f48f2d08eb4cf8b110",
X"4aaf6de5c79a0fe6c7f496d508e5e2f8b536",
X"4a06c2e5e3ba0fd9c3f49ee908e023f8b9a2",
X"495da8e600b60fcc2cf4a76808da0ef8be54",
X"48b422e61e8c0fbe05f4b05308d3a5f8c34c",
X"480a36e63d3b0faf4df4b9a808cce8f8c88a",
X"475fe6e65cc10fa007f4c36708c5d7f8ce0d",
X"46b535e67d1a0f9032f4cd9008be72f8d3d4",
X"460a28e69e460f7fd0f4d82108b6bbf8d9e1",
X"455ec3e6c0410f6ee3f4e31a08aeb1f8e032",
X"44b308e6e3090f5d6af4ee7b08a654f8e6c7",
X"4406fce7069d0f4b68f4fa42089da7f8ed9f",
X"435aa2e72af90f38ddf506700894a8f8f4bb",
X"42adffe7501d0f25caf51303088b58f8fc1a",
X"420115e776050f1230f51ffa0881b8f903bb",
X"4153e8e79cae0efe11f52d560877c8f90b9e",
X"40a67de7c4180ee96ef53b15086d89f913c4",
X"3ff8d6e7ec3f0ed448f549360862fcf91c2a",
X"3f4af8e815210ebea0f557ba085820f924d2",
X"3e9ce5e83ebc0ea877f5669e084cf7f92dba",
X"3deea3e8690d0e91cef575e3084181f936e2",
X"3d4034e894120e7aa8f585870835bef9404a",
X"3c919de8bfc90e6304f595890829b0f949f1",
X"3be2e0e8ec2f0e4ae5f5a5ea081d56f953d7",
X"3b3402e919420e324bf5b6a70810b2f95dfb",
X"3a8506e946ff0e1937f5c7c10803c3f9685d",
X"39d5f0e975640dffacf5d93607f68bf972fc",
X"3926c4e9a46e0de5aaf5eb0607e90af97dd8",
X"387785e9d41c0dcb33f5fd2f07db41f988f1",
X"37c837ea046a0db048f60fb107cd31f99445",
X"3718ddea35560d94ebf6228b07bed9f99fd5",
X"36697cea66dd0d791cf635bc07b03cf9ab9f",
X"35ba17ea98fe0d5cddf6494307a158f9b7a4",
X"350ab1eacbb50d4030f65d1f079230f9c3e2",
X"345b4eeaff000d2315f6714f0782c4f9d05a",
X"33abf3eb32dd0d058ff685d2077314f9dd0a",
X"32fca1eb67490ce79ff69aa8076322f9e9f2",
X"324d5eeb9c410cc945f6afcf0752edf9f712",
X"319e2debd1c30caa85f6c546074278fa0469",
X"30ef10ec07cd0c8b5ef6db0d0731c1fa11f6",
X"30400dec3e5b0c6bd3f6f1220720cbfa1fb8",
X"2f9126ec756c0c4be5f70784070f96fa2db0",
X"2ee25fecacfc0c2b95f71e3306fe22fa3bdc",
X"2e33bcece5090c0ae6f7352d06ec71fa4a3c",
X"2d8540ed1d910be9d7f74c7206da83fa58d0",
X"2cd6eeed56910bc86cf763ff06c859fa6796",
X"2c28cbed90060ba6a5f77bd506b5f4fa768e",
X"2b7adaedc9ee0b8484f793f206a355fa85b8",
X"2acd1eee04460b620bf7ac5506907cfa9512",
X"2a1f9aee3f0c0b3f3bf7c4fd067d6afaa49c",
X"297253ee7a3d0b1c15f7dde9066a20fab456",
X"28c54ceeb5d60af89cf7f7180656a0fac43f",
X"281888eef1d40ad4d0f810890642e8fad455",
X"276c0bef2e360ab0b4f82a3a062efcfae499",
X"26bfd8ef6af90a8c49f8442b061adbfaf50a",
X"2613f2efa8190a6790f85e5a060686fb05a7",
X"25685defe5950a428bf878c605f1fefb166f",
X"24bd1df0236a0a1d3cf8936f05dd45fb2761",
X"241234f0619409f7a4f8ae5305c85afb387e",
X"2367a7f0a01209d1c6f8c97005b33ffb49c4",
X"22bd78f0dee109aba2f8e4c7059df4fb5b32",
X"2213abf11dfe09853af9005505887bfb6cc8",
X"216a43f15d67095e8ff91c190572d5fb7e85",
X"20c144f19d190937a5f93813055d01fb9068",
X"2018b0f1dd1109107bf95440054702fba271",
X"1f708bf21d4d08e914f970a10530d9fbb49f",
X"1ec8d9f25dca08c171f98d33051a85fbc6f1",
X"1e219cf29e85089995f9a9f6050408fbd966",
X"1d7ad8f2df7d087180f9c6e804ed63fbebfe",
X"1cd48ff320ae084934f9e40904d697fbfeb7",
X"1c2ec6f362160820b4fa015604bfa5fc1192",
X"1b897ff3a3b207f800fa1ecf04a88dfc248d",
X"1ae4bef3e57f07cf1bfa3c72049151fc37a7",
X"1a4085f4277c07a605fa5a3f0479f2fc4ae0",
X"199cd8f469a4077cc1fa7834046270fc5e37",
X"18f9b9f4abf7075351fa9650044acdfc71ac",
X"18572df4ee710729b6fab492043309fc853c",
X"17b535f5310f06fff1fad2f7041b26fc98e9",
X"1713d6f573d006d605faf181040323fcacb0",
X"167311f5b6b006abf3fb102c03eb04fcc091",
X"15d2eaf5f9ad0681bcfb2ef803d2c7fcd48c",
X"153364f63cc5065763fb4de303ba6ffce89e",
X"149482f67ff5062ce9fb6ced03a1fcfcfcc9",
X"13f646f6c33a060251fb8c13038970fd110a",
X"1358b4f7069105d79afbab560370cafd2562",
X"12bbcff749f905acc8fbcab303580dfd39ce",
X"121f99f78d6f0581dbfbea29033f39fd4e4f",
X"118415f7d0f10556d7fc09b703264ffd62e4",
X"10e946f8147b052bbbfc295d030d50fd778b",
X"104f2ff8580b05008afc491702f43efd8c44",
X"0fb5d3f89b9f04d546fc68e602db18fda10f",
X"0f1d33f8df3504a9f1fc88c802c1e1fdb5ea",
X"0e8554f922c9047e8bfca8bc02a899fdcad4",
X"0dee38f9665b045317fcc8c1028f40fddfcd",
X"0d57e0f9a9e6042796fce8d40275d9fdf4d4",
X"0cc251f9ed6803fc0afd08f6025c64fe09e8",
X"0c2d8cfa30e003d074fd29250242e2fe1f08",
X"0b9994fa744b03a4d8fd495f022955fe3433",
X"0b066cfab7a6037934fd69a3020fbcfe4969",
X"0a7417fafaef034d8dfd89f101f619fe5ea9",
X"09e296fb3e240321e3fdaa4601dc6efe73f2",
X"0951ecfb814202f638fdcaa201c2bafe8943",
X"08c21cfbc44702ca8dfdeb0301a8fffe9e9b",
X"083328fc0730029ee5fe0b69018f3ffeb3f9",
X"07a512fc49fc027340fe2bd101757afec95d",
X"0717ddfc8ca80247a1fe4c3a015bb0fedec6",
X"068b8cfccf31021c09fe6ca50141e4fef433",
X"060020fd119601f079fe8d0e012815ff09a3",
X"05759cfd53d401c4f4fead75010e46ff1f15",
X"04ec01fd95e801997bfecdd900f477ff3489",
X"046353fdd7d2016e10feee3800daa8ff49fd",
X"03db94fe198d0142b3ff0e9200c0dcff5f71",
X"0354c5fe5b19011767ff2ee500a712ff74e4",
X"02cee9fe9c7300ec2eff4f2f008d4dff8a56",
X"024a02fedd9800c109ff6f7000738cff9fc4",
X"01c612ff1e870095f9ff8fa70059d1ffb530",
X"01431bff5f3d006b00ffafd100401dffca97",
X"00c11fff9fb900401fffcfef002671ffdff8",
X"004020ffdff8001559ffeffe000ccefff554");
	signal addr11,addr21: unsigned(7 downto 0);
begin
	addr11 <= addr1 when rising_edge(clk1);
	addr21 <= addr2 when rising_edge(clk2);
	q1 <= rom1(to_integer(addr11));
	q2 <= rom1(to_integer(addr21));
end architecture;
