library ieee;
library work;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
USE ieee.math_real.log2;
USE ieee.math_real.ceil;
use work.fft_types.all;

-- values are normalized to sqrt(n)
entity fft4_noPipeline is
	generic(dataBits: integer := 18);
	port(din: in complexArray(3 downto 0);
		dout: out complexArray(3 downto 0)
		);
end entity;

architecture a of fft4_noPipeline is
	signal a,b: complexArray(3 downto 0);
	signal resA1, resA2, resB1, resB2: complex;
	constant mask: integer := to_integer(signed'(dataBits-1 downto 0=>'1'));
begin
	a <= din;
	resA1 <= a(0) + a(2);
	resA2 <= a(0) - a(2);
	resB1 <= a(1) + a(3);
	resB2.re <= a(1).im - a(3).im;
	resB2.im <= a(3).re - a(1).re;
	
	b(0) <= resA1 + resB1;
	b(3) <= resA2 + resB2;
	b(2) <= resA1 - resB1;
	b(1) <= resA2 - resB2;
	
g:	for I in 0 to 3 generate
		dout(I) <= keepNBits(shift_right(b(I),1), dataBits);
	end generate;
end a;
