library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

--delay: 2 cycles
entity dsssCode1 is
	port(clk: in std_logic;
		addr: in unsigned(9 downto 0);
		data: out std_logic);
end entity;

architecture a of dsssCode1 is
	signal rom: std_logic_vector(1023 downto 0);
	signal addr1: unsigned(9 downto 0);
	signal data1: std_logic;
begin
	addr1 <= addr when rising_edge(clk);
	data1 <= rom(to_integer(addr1));
	data <= data1 when rising_edge(clk);
	rom <=
		"1000110000101011110011101001110110100011010010101011101111010001" &
		"1101110001111111001001001110100011011001101111110110110011110101" &
		"1111000010000111100000000001101100111000111110010100100101110001" &
		"0111010010010101100000000111000101011100000011001000010110111111" &
		"1000000010100011010001110000100000011111000110111010000110010011" &
		"1100000101011110011011111101101101010100011000010000111011100000" &
		"0010111110010010100101011101100111000000010101000010011110010100" &
		"0000000001010001010100101110111111101000101100100110100100001001" &
		"0100111000001001010011101111100110100000001110011010110001111010" &
		"1100010010110100011001000000010000101011101100111010011110101101" &
		"0010011011010010001100111101110000101010100001110000110100101010" &
		"0000101100011101010000001000101110011011011101011101100001010010" &
		"1010011001001111010011011001010111111100001000001111111101111101" &
		"0110100110011110011010110111110011010111001101001010011101010000" &
		"1101111101011011100110001111011111110101011110100100001110001001" &
		"1000111011101011110110101110010001110010001101000101111110000011";
end architecture;
