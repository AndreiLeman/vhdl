library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity usbtest2 is
    Port ( clk : in  STD_LOGIC);
end usbtest2;

architecture a of usbtest2 is

begin


end a;

